module UIDisplay();

endmodule