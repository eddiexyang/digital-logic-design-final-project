module VGADisplay

endmodule