module TopLevelShell();

endmodule