module KeyboardControl();

endmodule