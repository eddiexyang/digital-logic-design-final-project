module TopLevelShell();


endmodule