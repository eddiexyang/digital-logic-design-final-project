module FailureCheck(
    input [199:0] objects,
    input EN, // High-active enable signal
    output failure // 1 for failure, 0 for no failure
);

    genvar i, j;
    generate
        // TODO
    endgenerate
    integer i, j;
    
    clkdiv div_inst()


endmodule