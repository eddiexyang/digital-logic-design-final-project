module GameControl();

endmodule